LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY WH4574_OVERALL IS
	PORT(INVCC,S_H,S_M,S_S,CLK_5HZ,CLK1K : IN STD_LOGIC;
					LED_S0,LED_S1,LED_S2 : OUT STD_LOGIC;
		LED0,LED1,LED2,LED3,LED4,LED5,LED6,LED7 : OUT STD_LOGIC);
END WH4574_OVERALL;

ARCHITECTURE BEHAV OF WH4574_OVERALL IS
	COMPONENT WH4574_DIV5
		PORT(INCLK : IN STD_LOGIC;
				 Q : OUT STD_LOGIC);
	END COMPONENT;
	COMPONENT WH4574_DISPLAY
		PORT(DIN0,DIN1,DIN2,DIN3,DIN4,DIN5 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			CLK : IN STD_LOGIC;
			LED_SA,LED_SB,LED_SC : OUT STD_LOGIC;
			LED_A,LED_B,LED_C,LED_D,LED_E,LED_F,LED_G,LED_DP : OUT STD_LOGIC);
	END COMPONENT;
	COMPONENT WH4574_MUX2
		PORT(SEL,A,B :IN STD_LOGIC;
				Q : OUT STD_LOGIC);
	END COMPONENT;
	COMPONENT WH4574_COUNT60
		PORT(CLK : IN STD_LOGIC;
			BCD10,BCD1 : BUFFER STD_LOGIC_VECTOR(3 DOWNTO 0);
			PRESET : IN STD_LOGIC;
			CO : OUT STD_LOGIC);
	END COMPONENT;
	COMPONENT WH4574_COUNT24
		PORT(CLK : IN STD_LOGIC;
			BCD10,BCD1 : BUFFER STD_LOGIC_VECTOR(3 DOWNTO 0));
	END COMPONENT;
	COMPONENT WH4574_DIV40
		PORT(CLK : IN STD_LOGIC;
			  Q  : OUT STD_LOGIC);
	END COMPONENT;
	
	SIGNAL Q1,Q2,Q3,CO_S,CO_M : STD_LOGIC;
	SIGNAL H10,H1,M10,M1,S10,S1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
	
	BEGIN
	INST1:WH4574_MUX2 PORT MAP(SEL=>S_H,A=>CLK_5HZ,B=>CO_M,Q=>Q1);
	INST2:WH4574_MUX2 PORT MAP(SEL=>S_M,A=>CLK_5HZ,B=>CO_S,Q=>Q2);
	INST3:WH4574_DIV5 PORT MAP(INCLK=>CLK_5HZ,Q=>Q3);
	INST_H:WH4574_COUNT24 PORT MAP(CLK=>Q1,BCD10=>H10,BCD1=>H1);
	INST_M:WH4574_COUNT60 PORT MAP(CLK=>Q2,PRESET=>INVCC,BCD10=>M10,bcd1=>M1,CO=>CO_M);
	INST_S:WH4574_COUNT60 PORT MAP(CLK=>Q3,PRESET=>S_S,BCD10=>S10,bcd1=>S1,CO=>CO_S);
	INST_DISP:WH4574_DISPLAY PORT MAP(DIN5=>H10,DIN4=>H1,DIN3=>M10,DIN2=>M1,DIN1=>S10,DIN0=>S1,CLK=>CLK1K,
                                     LED_SA=>LED_S0,LED_SB=>LED_S1,LED_SC=>LED_S2,
                                     LED_A=>LED0,LED_B=>LED1,LED_C=>LED2,LED_D=>LED3,
                                     LED_E=>LED4,LED_F=>LED5,LED_G=>LED6,LED_DP=>LED7);
END ARCHITECTURE BEHAV;