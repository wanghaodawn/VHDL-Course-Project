LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY WH4574_COUNT60 IS
	PORT(
			CLK : IN STD_LOGIC;
			BCD10,BCD1 : BUFFER STD_LOGIC_VECTOR(3 DOWNTO 0);
			PRESET : IN STD_LOGIC;
			CO : OUT STD_LOGIC);
END WH4574_COUNT60;
ARCHITECTURE RTL OF WH4574_COUNT60 IS
	SIGNAL CO_1 : STD_LOGIC;
	BEGIN
		PROCESS(CLK,PRESET)
		BEGIN
			IF PRESET = '0' THEN
				BCD1 <= "0000";
			ELSE
				IF CLK = '1' AND CLK'EVENT THEN
					IF BCD1 = "1001" THEN
						BCD1 <= "0000";
					ELSE
					BCD1 <= BCD1 + 1;
					END IF;
				END IF;
			END IF;
		END PROCESS;
		
		PROCESS(CLK,PRESET,BCD1)
		BEGIN
			IF PRESET = '0' THEN
				BCD10 <= "0000";
				CO_1 <= '0';
			ELSE
				IF CLK = '1' AND CLK'EVENT THEN
					IF BCD1 = "1000" AND BCD10 = "0101" THEN
						CO_1 <= '1';
					ELSIF BCD1 = "1001" AND BCD10 = "0101" THEN
						BCD10 <= "0000";
						CO_1 <= '0';
					ELSIF BCD1 = "1001" THEN
						BCD10 <= BCD10 + '1';
						CO_1 <= '0';
					END IF;
				END IF;
			END IF;
		END PROCESS;
		
		CO <= NOT CO_1;
		
		END RTL;
						