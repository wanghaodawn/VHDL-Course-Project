LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY WH4574_DISPLAY IS
 PORT(DIN0,DIN1,DIN2,DIN3,DIN4,DIN5 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      CLK : IN STD_LOGIC;
      LED_SA,LED_SB,LED_SC : OUT STD_LOGIC;
      LED_A,LED_B,LED_C,LED_D,LED_E,LED_F,LED_G,LED_DP : OUT STD_LOGIC);
  END ENTITY WH4574_DISPLAY;

ARCHITECTURE behav of WH4574_DISPLAY IS
	SIGNAL SEG : STD_LOGIC_VECTOR(6 DOWNTO 0); 
	SIGNAL SEL : STD_LOGIC_VECTOR(2 DOWNTO 0);
	SIGNAL NUM : STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL S   : STD_LOGIC_VECTOR(2 DOWNTO 0);
  
   BEGIN
    LED_SA <= SEL(0);
    LED_SB <= SEL(1);
    LED_SC <= SEL(2);
    LED_A <= SEG(0);
    LED_B <= SEG(1);
    LED_C <= SEG(2);
    LED_D <= SEG(3);
    LED_E <= SEG(4);
    LED_F <= SEG(5);
    LED_G <= SEG(6);
  
	PROCESS(CLK)
	BEGIN
		IF CLK'EVENT AND CLK = '1' THEN
			IF S = "101" THEN
				S <= "000";
			ELSE
				S <= S + '1';
			END IF;
		END IF;
	END PROCESS;
   
	PROCESS(S,DIN0,DIN1,DIN2,DIN3,DIN4,DIN5)
    BEGIN
		IF S = "000" THEN
			SEL <= "000";
            NUM <= DIN0;
            LED_DP <= '0';
			ELSIF S = "001" THEN
				SEL <= "001";
				NUM <= DIN1;
				LED_DP <= '0';
				ELSIF S = "010" THEN
					SEL <= "010";
					NUM <= DIN2;
					LED_DP <= '0';
					ELSIF S = "011" THEN
					SEL <= "011";
					NUM <= DIN3;
					LED_DP <= '0';
						ELSIF S="100" THEN
						SEL <= "100";
						NUM <= DIN4;
						LED_DP <= '0';
							ELSIF S = "101" THEN
								SEL <= "101";
								NUM <= DIN5;
								LED_DP <= '0';
								ELSE 
									SEL <= "XXX";
									NUM <= "XXXX";
									LED_DP <= '0';
		END IF;
	END PROCESS;
  
	SEG<="0111111" WHEN NUM = 0 ELSE
		"0000110" WHEN NUM = 1 ELSE
		"1011011" WHEN NUM = 2 ELSE
		"1001111" WHEN NUM = 3 ELSE
		"1100110" WHEN NUM = 4 ELSE
		"1101101" WHEN NUM = 5 ELSE
		"1111101" WHEN NUM = 6 ELSE
		"0000111" WHEN NUM = 7 ELSE
		"1111111" WHEN NUM = 8 ELSE
		"1101111" WHEN NUM = 9 ELSE
		"1110111" WHEN NUM = 10 ELSE
		"1111100" WHEN NUM = 11 ELSE
		"0111001" WHEN NUM = 12 ELSE
		"1011110" WHEN NUM = 13 ELSE
		"1111001" WHEN NUM = 14 ELSE
		"1110001" WHEN NUM = 15 ELSE
		"0000000";
END behav;