LIBRARY IEEE;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY WH4574_DIV4K IS
 PORT(CLK:IN STD_LOGIC;
      OUTCLK:OUT STD_LOGIC);
END ENTITY;
ARCHITECTURE BEHAV OF WH4574_DIV4K IS
 SIGNAL COUNT:INTEGER RANGE 0 TO 1999;
 SIGNAL Q1,COUNT2:STD_LOGIC;
  BEGIN
   PROCESS(CLK)
    BEGIN
    IF CLK'EVENT AND CLK='1' THEN
      IF COUNT=1999 THEN
         COUNT<=0;
         Q1<='1';
      ELSE 
       COUNT<=COUNT+1;
           Q1<='0';
       END IF;
    END IF;
   END PROCESS;
   PROCESS(Q1)
    BEGIN
     IF Q1'EVENT AND Q1='1' THEN
      COUNT2<=NOT COUNT2;
      END IF;
   END PROCESS;
   OUTCLK<=COUNT2;
   END BEHAV;