LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY WH4574_DIV4 IS
	PORT(
			CLK : IN STD_LOGIC;
			Q : OUT STD_LOGIC);
END WH4574_DIV4;
ARCHITECTURE RTL OF WH4574_DIV4 IS
	SIGNAL CC : INTEGER RANGE 0 TO 3;
	BEGIN
		PROCESS(CLK)
		BEGIN
			IF CLK = '1' AND CLK'EVENT THEN
				CASE CC IS
					WHEN 0 => CC <= CC + 1;Q <= '0';
					WHEN 1 => CC <= CC + 1;Q <= '0';
					WHEN 2 => CC <= CC + 1;Q <= '1';
					WHEN 3 => CC <= 0;     Q <= '1';
				END CASE;
			END IF;
		END PROCESS;	
END RTL;
						