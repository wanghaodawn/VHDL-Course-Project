LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY WH4574_DIV5 IS
	PORT(INCLK : IN STD_LOGIC;
			 Q : OUT STD_LOGIC);
END ENTITY WH4574_DIV5;

ARCHITECTURE behav of WH4574_DIV5 IS
	SIGNAL COUNT : STD_LOGIC_VECTOR(2 DOWNTO 0);
	SIGNAL CLK, OUTCLK1, DIVIDE2, DIVIDE3, OUTCLK2 : STD_LOGIC;
	BEGIN
	CLK <= INCLK XOR DIVIDE2;
    PROCESS(CLK)
	BEGIN
		IF CLK'EVENT AND CLK = '1' THEN
			IF COUNT = "000" THEN
				COUNT <= "011"-1;
				OUTCLK1 <= '1';
			ELSE
				COUNT <= COUNT-1;
				OUTCLK1 <= '0';
			END IF;
		END IF;
    END PROCESS;
    
    PROCESS(OUTCLK1)
    BEGIN
		IF OUTCLK1'EVENT AND OUTCLK1 = '1' THEN
			DIVIDE2 <= NOT DIVIDE2;
        END IF;
    END PROCESS;
   
    Q <= DIVIDE2;  
    
END behav;    
     