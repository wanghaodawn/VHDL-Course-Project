LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY WH4574_DIV2 IS
	PORT(CLK : IN STD_LOGIC;
			 Q : OUT STD_LOGIC);
END ENTITY WH4574_DIV2;

ARCHITECTURE BEHAV OF WH4574_DIV2 IS
	SIGNAL COUNT : STD_LOGIC;
	SIGNAL QQ : STD_LOGIC;
	BEGIN

    PROCESS(CLK)
	BEGIN
		IF CLK'EVENT AND CLK = '1' THEN
				QQ <= NOT QQ;
		END IF;
    END PROCESS;
    
    Q <= QQ;
END BEHAV;    
     