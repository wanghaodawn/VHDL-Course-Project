LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY WH4574_SEL2 IS
	PORT(
			CLK : IN STD_LOGIC;
			SEL : IN STD_LOGIC;
			Q : OUT STD_LOGIC);
END WH4574_SEL2;
ARCHITECTURE RTL OF WH4574_SEL2 IS
	SIGNAL C : INTEGER RANGE 0 TO 50;
	BEGIN
		PROCESS(SEL,CLK)
		BEGIN
		IF SEL = '0' THEN
			Q <= CLK;
		ELSE
			IF CLK'EVENT AND CLK = '1' THEN
				IF C = 50 THEN
					Q <= CLK;
					C <= 0;
				ELSE
					C <= C + 1;
					Q <= '1';
				END IF;
			END IF;
		END IF;
		END PROCESS;	
END RTL;
						