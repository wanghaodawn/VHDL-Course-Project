LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY WH4574_KEYIN IS
	PORT(CLK,KEY : IN STD_LOGIC;
			 Q : OUT STD_LOGIC);
END ENTITY WH4574_KEYIN;

ARCHITECTURE BEHAV OF WH4574_KEYIN IS
	SIGNAL COUNT : INTEGER RANGE 0 TO 2;
	BEGIN

    PROCESS(CLK)
	BEGIN
		IF CLK'EVENT AND CLK = '1' THEN
			CASE COUNT IS
				WHEN 0 => IF KEY = '0' THEN
							COUNT <= 1;
							Q <= '1';
						  END IF;
				WHEN 1 => IF KEY = '0' THEN
							COUNT <= 2;
							Q <= '0';
						  END IF;
				WHEN 2 => IF KEY = '1' THEN
							COUNT <= 0;
							Q <= '1';
						  END IF;
			END CASE;
		END IF;
	END PROCESS;
END BEHAV;    
     