LIBRARY IEEE;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY WH4574_DIV2K_CTRL IS
 PORT(Q_1K,Q_2K,CLK50M:IN STD_LOGIC;
      CLK_BEEP:OUT STD_LOGIC);
END ENTITY;
ARCHITECTURE BEHAV OF WH4574_DIV2K_CTRL IS
 SIGNAL COUNT1:INTEGER RANGE 0 TO 2499;
 SIGNAL COUNT2:STD_LOGIC; 
 SIGNAL CO:STD_LOGIC; 
       BEGIN
  PROCESS(CLK50M)
   BEGIN
   IF CLK50M'EVENT AND CLK50M='1' THEN
    IF Q_2K = '1' THEN
    	IF COUNT1=1249 THEN
		COUNT1<=0;
		CO<='1';
		ELSE 
		COUNT1<=COUNT1+1;
		CO<='0';
		END IF;
    ELSIF Q_1K = '1' THEN
		IF COUNT1=2499 THEN
		COUNT1<=0;
		CO<='1';
		ELSE 
		COUNT1<=COUNT1+1;
		CO<='0';
		END IF;
   END IF;
   END IF;
  END PROCESS;
   PROCESS(CO)
     BEGIN
     IF CO'EVENT AND CO='1' THEN
      COUNT2<=NOT COUNT2;
     END IF;
   END PROCESS;
   CLK_BEEP<=COUNT2;
END BEHAV;